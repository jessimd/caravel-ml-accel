magic
tech sky130B
magscale 1 2
timestamp 1660091864
<< obsli1 >>
rect 1104 2159 398820 597329
<< obsm1 >>
rect 14 2128 399726 597360
<< metal2 >>
rect 2594 599200 2650 600000
rect 27710 599200 27766 600000
rect 52182 599200 52238 600000
rect 77298 599200 77354 600000
rect 101770 599200 101826 600000
rect 126886 599200 126942 600000
rect 152002 599200 152058 600000
rect 176474 599200 176530 600000
rect 201590 599200 201646 600000
rect 226062 599200 226118 600000
rect 251178 599200 251234 600000
rect 276294 599200 276350 600000
rect 300766 599200 300822 600000
rect 325882 599200 325938 600000
rect 350354 599200 350410 600000
rect 375470 599200 375526 600000
rect 399942 599200 399998 600000
rect 18 0 74 800
rect 24490 0 24546 800
rect 49606 0 49662 800
rect 74078 0 74134 800
rect 99194 0 99250 800
rect 123666 0 123722 800
rect 148782 0 148838 800
rect 173898 0 173954 800
rect 198370 0 198426 800
rect 223486 0 223542 800
rect 247958 0 248014 800
rect 273074 0 273130 800
rect 298190 0 298246 800
rect 322662 0 322718 800
rect 347778 0 347834 800
rect 372250 0 372306 800
rect 397366 0 397422 800
<< obsm2 >>
rect 20 599144 2538 599298
rect 2706 599144 27654 599298
rect 27822 599144 52126 599298
rect 52294 599144 77242 599298
rect 77410 599144 101714 599298
rect 101882 599144 126830 599298
rect 126998 599144 151946 599298
rect 152114 599144 176418 599298
rect 176586 599144 201534 599298
rect 201702 599144 226006 599298
rect 226174 599144 251122 599298
rect 251290 599144 276238 599298
rect 276406 599144 300710 599298
rect 300878 599144 325826 599298
rect 325994 599144 350298 599298
rect 350466 599144 375414 599298
rect 375582 599144 399886 599298
rect 20 856 399942 599144
rect 130 800 24434 856
rect 24602 800 49550 856
rect 49718 800 74022 856
rect 74190 800 99138 856
rect 99306 800 123610 856
rect 123778 800 148726 856
rect 148894 800 173842 856
rect 174010 800 198314 856
rect 198482 800 223430 856
rect 223598 800 247902 856
rect 248070 800 273018 856
rect 273186 800 298134 856
rect 298302 800 322606 856
rect 322774 800 347722 856
rect 347890 800 372194 856
rect 372362 800 397310 856
rect 397478 800 399942 856
<< metal3 >>
rect 0 576648 800 576768
rect 399200 573928 400000 574048
rect 0 550808 800 550928
rect 399200 547408 400000 547528
rect 0 524288 800 524408
rect 399200 521568 400000 521688
rect 0 498448 800 498568
rect 399200 495048 400000 495168
rect 0 471928 800 472048
rect 399200 469208 400000 469328
rect 0 446088 800 446208
rect 399200 442688 400000 442808
rect 0 419568 800 419688
rect 399200 416168 400000 416288
rect 0 393048 800 393168
rect 399200 390328 400000 390448
rect 0 367208 800 367328
rect 399200 363808 400000 363928
rect 0 340688 800 340808
rect 399200 337968 400000 338088
rect 0 314848 800 314968
rect 399200 311448 400000 311568
rect 0 288328 800 288448
rect 399200 284928 400000 285048
rect 0 261808 800 261928
rect 399200 259088 400000 259208
rect 0 235968 800 236088
rect 399200 232568 400000 232688
rect 0 209448 800 209568
rect 399200 206728 400000 206848
rect 0 183608 800 183728
rect 399200 180208 400000 180328
rect 0 157088 800 157208
rect 399200 153688 400000 153808
rect 0 130568 800 130688
rect 399200 127848 400000 127968
rect 0 104728 800 104848
rect 399200 101328 400000 101448
rect 0 78208 800 78328
rect 399200 75488 400000 75608
rect 0 52368 800 52488
rect 399200 48968 400000 49088
rect 0 25848 800 25968
rect 399200 23128 400000 23248
<< obsm3 >>
rect 800 576848 399200 597345
rect 880 576568 399200 576848
rect 800 574128 399200 576568
rect 800 573848 399120 574128
rect 800 551008 399200 573848
rect 880 550728 399200 551008
rect 800 547608 399200 550728
rect 800 547328 399120 547608
rect 800 524488 399200 547328
rect 880 524208 399200 524488
rect 800 521768 399200 524208
rect 800 521488 399120 521768
rect 800 498648 399200 521488
rect 880 498368 399200 498648
rect 800 495248 399200 498368
rect 800 494968 399120 495248
rect 800 472128 399200 494968
rect 880 471848 399200 472128
rect 800 469408 399200 471848
rect 800 469128 399120 469408
rect 800 446288 399200 469128
rect 880 446008 399200 446288
rect 800 442888 399200 446008
rect 800 442608 399120 442888
rect 800 419768 399200 442608
rect 880 419488 399200 419768
rect 800 416368 399200 419488
rect 800 416088 399120 416368
rect 800 393248 399200 416088
rect 880 392968 399200 393248
rect 800 390528 399200 392968
rect 800 390248 399120 390528
rect 800 367408 399200 390248
rect 880 367128 399200 367408
rect 800 364008 399200 367128
rect 800 363728 399120 364008
rect 800 340888 399200 363728
rect 880 340608 399200 340888
rect 800 338168 399200 340608
rect 800 337888 399120 338168
rect 800 315048 399200 337888
rect 880 314768 399200 315048
rect 800 311648 399200 314768
rect 800 311368 399120 311648
rect 800 288528 399200 311368
rect 880 288248 399200 288528
rect 800 285128 399200 288248
rect 800 284848 399120 285128
rect 800 262008 399200 284848
rect 880 261728 399200 262008
rect 800 259288 399200 261728
rect 800 259008 399120 259288
rect 800 236168 399200 259008
rect 880 235888 399200 236168
rect 800 232768 399200 235888
rect 800 232488 399120 232768
rect 800 209648 399200 232488
rect 880 209368 399200 209648
rect 800 206928 399200 209368
rect 800 206648 399120 206928
rect 800 183808 399200 206648
rect 880 183528 399200 183808
rect 800 180408 399200 183528
rect 800 180128 399120 180408
rect 800 157288 399200 180128
rect 880 157008 399200 157288
rect 800 153888 399200 157008
rect 800 153608 399120 153888
rect 800 130768 399200 153608
rect 880 130488 399200 130768
rect 800 128048 399200 130488
rect 800 127768 399120 128048
rect 800 104928 399200 127768
rect 880 104648 399200 104928
rect 800 101528 399200 104648
rect 800 101248 399120 101528
rect 800 78408 399200 101248
rect 880 78128 399200 78408
rect 800 75688 399200 78128
rect 800 75408 399120 75688
rect 800 52568 399200 75408
rect 880 52288 399200 52568
rect 800 49168 399200 52288
rect 800 48888 399120 49168
rect 800 26048 399200 48888
rect 880 25768 399200 26048
rect 800 23328 399200 25768
rect 800 23048 399120 23328
rect 800 2143 399200 23048
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
rect 50288 2128 50608 597360
rect 65648 2128 65968 597360
rect 81008 2128 81328 597360
rect 96368 2128 96688 597360
rect 111728 2128 112048 597360
rect 127088 2128 127408 597360
rect 142448 2128 142768 597360
rect 157808 2128 158128 597360
rect 173168 2128 173488 597360
rect 188528 2128 188848 597360
rect 203888 2128 204208 597360
rect 219248 2128 219568 597360
rect 234608 2128 234928 597360
rect 249968 2128 250288 597360
rect 265328 2128 265648 597360
rect 280688 2128 281008 597360
rect 296048 2128 296368 597360
rect 311408 2128 311728 597360
rect 326768 2128 327088 597360
rect 342128 2128 342448 597360
rect 357488 2128 357808 597360
rect 372848 2128 373168 597360
rect 388208 2128 388528 597360
<< obsm4 >>
rect 83779 2347 96288 597005
rect 96768 2347 111648 597005
rect 112128 2347 127008 597005
rect 127488 2347 142368 597005
rect 142848 2347 157728 597005
rect 158208 2347 173088 597005
rect 173568 2347 188448 597005
rect 188928 2347 203808 597005
rect 204288 2347 219168 597005
rect 219648 2347 234528 597005
rect 235008 2347 249888 597005
rect 250368 2347 265248 597005
rect 265728 2347 280608 597005
rect 281088 2347 295968 597005
rect 296448 2347 306485 597005
<< labels >>
rlabel metal3 s 0 261808 800 261928 6 clock_clock
port 1 nsew signal input
rlabel metal2 s 201590 599200 201646 600000 6 custom_boot
port 2 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 jtag_TCK
port 3 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 jtag_TDI
port 4 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 jtag_TDO
port 5 nsew signal output
rlabel metal3 s 399200 469208 400000 469328 6 jtag_TMS
port 6 nsew signal input
rlabel metal2 s 372250 0 372306 800 6 reset
port 7 nsew signal input
rlabel metal3 s 399200 521568 400000 521688 6 serial_tl_bits_in_bits[0]
port 8 nsew signal input
rlabel metal3 s 399200 232568 400000 232688 6 serial_tl_bits_in_bits[10]
port 9 nsew signal input
rlabel metal3 s 0 524288 800 524408 6 serial_tl_bits_in_bits[11]
port 10 nsew signal input
rlabel metal3 s 399200 23128 400000 23248 6 serial_tl_bits_in_bits[12]
port 11 nsew signal input
rlabel metal2 s 350354 599200 350410 600000 6 serial_tl_bits_in_bits[13]
port 12 nsew signal input
rlabel metal2 s 52182 599200 52238 600000 6 serial_tl_bits_in_bits[14]
port 13 nsew signal input
rlabel metal3 s 399200 75488 400000 75608 6 serial_tl_bits_in_bits[15]
port 14 nsew signal input
rlabel metal3 s 0 314848 800 314968 6 serial_tl_bits_in_bits[16]
port 15 nsew signal input
rlabel metal3 s 399200 311448 400000 311568 6 serial_tl_bits_in_bits[17]
port 16 nsew signal input
rlabel metal3 s 399200 390328 400000 390448 6 serial_tl_bits_in_bits[18]
port 17 nsew signal input
rlabel metal3 s 0 288328 800 288448 6 serial_tl_bits_in_bits[19]
port 18 nsew signal input
rlabel metal3 s 399200 259088 400000 259208 6 serial_tl_bits_in_bits[1]
port 19 nsew signal input
rlabel metal2 s 375470 599200 375526 600000 6 serial_tl_bits_in_bits[20]
port 20 nsew signal input
rlabel metal3 s 399200 206728 400000 206848 6 serial_tl_bits_in_bits[21]
port 21 nsew signal input
rlabel metal2 s 226062 599200 226118 600000 6 serial_tl_bits_in_bits[22]
port 22 nsew signal input
rlabel metal3 s 399200 153688 400000 153808 6 serial_tl_bits_in_bits[23]
port 23 nsew signal input
rlabel metal2 s 298190 0 298246 800 6 serial_tl_bits_in_bits[24]
port 24 nsew signal input
rlabel metal3 s 399200 442688 400000 442808 6 serial_tl_bits_in_bits[25]
port 25 nsew signal input
rlabel metal3 s 399200 495048 400000 495168 6 serial_tl_bits_in_bits[26]
port 26 nsew signal input
rlabel metal2 s 397366 0 397422 800 6 serial_tl_bits_in_bits[27]
port 27 nsew signal input
rlabel metal3 s 0 419568 800 419688 6 serial_tl_bits_in_bits[28]
port 28 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 serial_tl_bits_in_bits[29]
port 29 nsew signal input
rlabel metal2 s 251178 599200 251234 600000 6 serial_tl_bits_in_bits[2]
port 30 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 serial_tl_bits_in_bits[30]
port 31 nsew signal input
rlabel metal3 s 0 393048 800 393168 6 serial_tl_bits_in_bits[31]
port 32 nsew signal input
rlabel metal3 s 399200 416168 400000 416288 6 serial_tl_bits_in_bits[3]
port 33 nsew signal input
rlabel metal2 s 77298 599200 77354 600000 6 serial_tl_bits_in_bits[4]
port 34 nsew signal input
rlabel metal3 s 0 550808 800 550928 6 serial_tl_bits_in_bits[5]
port 35 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 serial_tl_bits_in_bits[6]
port 36 nsew signal input
rlabel metal2 s 347778 0 347834 800 6 serial_tl_bits_in_bits[7]
port 37 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 serial_tl_bits_in_bits[8]
port 38 nsew signal input
rlabel metal3 s 399200 101328 400000 101448 6 serial_tl_bits_in_bits[9]
port 39 nsew signal input
rlabel metal2 s 101770 599200 101826 600000 6 serial_tl_bits_in_ready
port 40 nsew signal output
rlabel metal3 s 0 498448 800 498568 6 serial_tl_bits_in_valid
port 41 nsew signal input
rlabel metal3 s 399200 48968 400000 49088 6 serial_tl_bits_out_bits[0]
port 42 nsew signal output
rlabel metal2 s 126886 599200 126942 600000 6 serial_tl_bits_out_bits[10]
port 43 nsew signal output
rlabel metal3 s 399200 180208 400000 180328 6 serial_tl_bits_out_bits[11]
port 44 nsew signal output
rlabel metal3 s 399200 284928 400000 285048 6 serial_tl_bits_out_bits[12]
port 45 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 serial_tl_bits_out_bits[13]
port 46 nsew signal output
rlabel metal3 s 0 367208 800 367328 6 serial_tl_bits_out_bits[14]
port 47 nsew signal output
rlabel metal3 s 0 471928 800 472048 6 serial_tl_bits_out_bits[15]
port 48 nsew signal output
rlabel metal2 s 176474 599200 176530 600000 6 serial_tl_bits_out_bits[16]
port 49 nsew signal output
rlabel metal2 s 223486 0 223542 800 6 serial_tl_bits_out_bits[17]
port 50 nsew signal output
rlabel metal2 s 18 0 74 800 6 serial_tl_bits_out_bits[18]
port 51 nsew signal output
rlabel metal2 s 273074 0 273130 800 6 serial_tl_bits_out_bits[19]
port 52 nsew signal output
rlabel metal2 s 152002 599200 152058 600000 6 serial_tl_bits_out_bits[1]
port 53 nsew signal output
rlabel metal2 s 276294 599200 276350 600000 6 serial_tl_bits_out_bits[20]
port 54 nsew signal output
rlabel metal2 s 399942 599200 399998 600000 6 serial_tl_bits_out_bits[21]
port 55 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 serial_tl_bits_out_bits[22]
port 56 nsew signal output
rlabel metal3 s 0 340688 800 340808 6 serial_tl_bits_out_bits[23]
port 57 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 serial_tl_bits_out_bits[24]
port 58 nsew signal output
rlabel metal3 s 399200 573928 400000 574048 6 serial_tl_bits_out_bits[25]
port 59 nsew signal output
rlabel metal3 s 0 209448 800 209568 6 serial_tl_bits_out_bits[26]
port 60 nsew signal output
rlabel metal2 s 198370 0 198426 800 6 serial_tl_bits_out_bits[27]
port 61 nsew signal output
rlabel metal3 s 399200 547408 400000 547528 6 serial_tl_bits_out_bits[28]
port 62 nsew signal output
rlabel metal3 s 399200 127848 400000 127968 6 serial_tl_bits_out_bits[29]
port 63 nsew signal output
rlabel metal2 s 2594 599200 2650 600000 6 serial_tl_bits_out_bits[2]
port 64 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 serial_tl_bits_out_bits[30]
port 65 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 serial_tl_bits_out_bits[31]
port 66 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 serial_tl_bits_out_bits[3]
port 67 nsew signal output
rlabel metal3 s 0 235968 800 236088 6 serial_tl_bits_out_bits[4]
port 68 nsew signal output
rlabel metal3 s 399200 363808 400000 363928 6 serial_tl_bits_out_bits[5]
port 69 nsew signal output
rlabel metal2 s 247958 0 248014 800 6 serial_tl_bits_out_bits[6]
port 70 nsew signal output
rlabel metal2 s 325882 599200 325938 600000 6 serial_tl_bits_out_bits[7]
port 71 nsew signal output
rlabel metal2 s 300766 599200 300822 600000 6 serial_tl_bits_out_bits[8]
port 72 nsew signal output
rlabel metal3 s 0 576648 800 576768 6 serial_tl_bits_out_bits[9]
port 73 nsew signal output
rlabel metal2 s 27710 599200 27766 600000 6 serial_tl_bits_out_ready
port 74 nsew signal input
rlabel metal2 s 322662 0 322718 800 6 serial_tl_bits_out_valid
port 75 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 serial_tl_clock
port 76 nsew signal output
rlabel metal3 s 0 446088 800 446208 6 uart_0_rxd
port 77 nsew signal input
rlabel metal3 s 399200 337968 400000 338088 6 uart_0_txd
port 78 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 597360 6 vccd1
port 79 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 597360 6 vssd1
port 80 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 597360 6 vssd1
port 80 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 400000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 203801980
string GDS_FILE /home/ubuntu/caravel-ml-accel/openlane/ChipTop/runs/22_08_09_23_16/results/signoff/ChipTop.magic.gds
string GDS_START 1642294
<< end >>

